SLVM023 (PSpice format)
**************************************
**  This file was created by TINA   **
**         www.tina.com             **
**      (c) DesignSoft, Inc.        **
**     www.designsoftware.com       **
**************************************
*.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\EXAMPLES\SPICE\TSPICE.LIB"
*.LIB "C:\Program Files (x86)\DesignSoft\Tina 9 - TI\SPICELIB\Operational Amplifiers.LIB"
.LIB tps40200p.lib
.TEMP 27
*.AC DEC 20 10 1MEG
.TRAN 1.4U 700U UIC

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=14
.PROBE V([N5R2V]) V([VISEN]) V([VSW]) V([VSTART]) V([VRC])
.PROBE V([VGATE])

VIN_12      8 0 12
XU1         VRC VSTART 3 4 N5R2V 6 VISEN 8 TPS40200
Rc108       9 N5R2V 2M
Rc107       10 N5R2V 2M
XT1         VSW VGATE 11 12 FDS4685_0
XD1         N5R2V VSW SS10P4_0
RL          0 N5R2V 2.08
R1          12 0 34K
C104        3 4 150P IC=0
C103        3 15 5.6N IC=0
C109        4 16 2.2N IC=0
R105        15 4 3.48K
R111        N5R2V 4 1.54K
R108        16 0 226
R109        4 0 10K
C105        VSTART N5R2V 18N IC=0
C108        VRC N5R2V 620P IC=0
R101        8 VRC 34K
C108_2      0 9 47U IC=0
C106        8 N5R2V 100N IC=0
C107        0 10 47U IC=0
R103        6 VGATE 2
R102        VISEN 11 1K
C100        8 VISEN 100P IC=0
R100        8 11 10M
C101        8 0 10U IC=0
L100        VSW 0 5.2U IC=1


* SUBCKT: TPS40200 encrypted macro, content not displayed


*FDS4685 AT TEMP. ELECTRICAL MODEL
*-----------------------------------------------------
.SUBCKT FDS4685_0  20 10 30 50
*20=DRAIN 10=GATE 30=SOURCE 50=VTEMP
RG 10 11X 1
RDU 12X 1 1U
M1 2 1 4X 4X DMOS L=1U W=1U
.MODEL DMOS PMOS(VTO=-1.7 KP=2.6E+1 THETA=.1 VMAX=5.5E5 LEVEL=3)
CGS 1 5X 1736P
RD 20 4 6E-3
DDS 4 5X DDS
.MODEL DDS D(M=5.1E-1 VJ=1.03E-1 CJO=570P)
DBODY 20 5X DBODY
.MODEL DBODY D(IS=2.86E-13 N=0.932967 RS=1.3E-4 TT=12.41N)
RA 4 2 6E-3
RS 5X 5 0.5M
LS 5 30 0.5N
M2 1 8 6 6 INTER
E2 8 6 4 1 2
.MODEL INTER PMOS(VTO=0 KP=10 LEVEL=1)
CGDMAX 7 4 1329P
RCGD 7 4 10MEG
DGD 4 6 DGD
RDGD 4 6 10MEG
.MODEL DGD D(M=2.69E-1 VJ=8.56E-3 CJO=1329P)
M3 7 9 1 1 INTER
E3 9 1 4 1 -2
*ZX SECTION
EOUT 4X 6X POLY(2) (1X,0) (3X,0) 0 0 0 0 1
FCOPY 0 3X VSENSE 1
RIN 1X 0 1G
VSENSE 6X 5X 0
RREF 3X 0 10M
*TEMP SECTION
ED 101 0 VALUE {V(50,100)}
VAMB 100 0 25
EKP 1X 0 101 0 .012
*VTO TEMP SECTION
EVTO 102 0 101 0 .005
EVT 11X 12X 102 0 1
*DIODE THEMO BREAKDOWN SECTION
EBL VB1 VB2 101 0 .08
VBLK VB2 0 40
D DB1 20 DBLK
.MODEL DBLK D(IS=1E-14 CJO=.1P RS=.1)
EDB 0 DB1 VB1 0 1
.ENDS FDS4685_0
*FDS4685 (REV.A) 8/25/05
*ST



**********************************
* COPYRIGHT:                     *
*   THOMATRONIK GMBH, GERMANY    *
*   INFO@THOMATRONIK.DE          *
**********************************
*   PSPICE
.SUBCKT SS10P4_0  A C
DDIO A C LEGD
DGR A C GRD
.MODEL LEGD D IS = 1.00002E-015 N = 0.663355 RS = 0.00362975
+ EG = 0.400729 XTI = 0.500158 T_MEASURED = 27
+ CJO = 2.15315E-009 VJ = 0.7 M = 0.539076 FC = 0.5
+ TT = 2.4663E-010 BV = 44 IBV = 0.1 AF = 1 KF = 0
.MODEL GRD D IS = 5.36639E-006 N = 0.947898 RS = 0.0132545
+ EG = 0.663278 XTI = 0.539193 T_MEASURED = 27
.ENDS



.END
