* Experiment 1: Opamp

* INPUT SIGNAL
VG vg 0 PULSE(0 1 1u 10n 10n 1u 2u 4)

* SUPPLY
VDD vdd 0 10
VSS 0 vss 10

XU1 vg vf1 vdd vss vf1 tl082
XU2 vg N001 vdd vss vf2 tl082
XU3 0 N002 vdd vss vf3 tl082

R1 N001 0 1k
R2 vf2 N001 2k
R3 N002 vg 1k
R4 vf3 N002 2k

* MODEL
.inc tl082.cir

* ANALYSIS
.tran 10u

.end
