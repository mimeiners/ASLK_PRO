AGC
**************************************
**  This file was created by TINA   **
**         www.tina.com             **
**      (c) DesignSoft, Inc.        **
**     www.designsoftware.com       **
**************************************


*.TEMP 27
*.AC DEC 20 10 1MEG
.TRAN 60U 30M
*.DC LIN V_Ref 0 1 10M

.save all


* Power Supply
VDD	        vdd 0 10
VSS         vss 0 -10
VE          ve  0 10

Vref        inp 0 DC 0
+                 SIN( 0 3 50 0 0 0 )

* Signals
Vin         vin 0 DC 0
+                 AC 1 0
+                 SIN( 0 5 50 0 0 0 )


* Multiplier 1
Xmult1      vin 0 ve vfb 0 vdd vo1 z11 0 vss MPY634_BEHAVIORAL_0
Rvo1        vo1 z11 90K
Rz11        z11 0   10K
Cz11        z11 0   200P

* Multiplier 2
Xmult2      vo1 0 ve vo1 0 vdd vo2 z12 0 vss MPY634_BEHAVIORAL_0
Rvo2        vo2 z12 90K
Rz12        z12 0   10K
Cz12        z12 0   200P

* Low pass
Rlp          vo3 vo2 1K
Clp          vo3 0   10U

* Comparator
Xcomp       inp vo3 vdd vss vo3 TL082_0



* TL082 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 06/16/89 AT 13:08
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* ------------------------------------------------------------------------
*|(C) COPYRIGHT TEXAS INSTRUMENTS INCORPORATED 2007. ALL RIGHTS RESERVED. |
*|                                                                        |
*|THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.    |
*|NO WARRANTIES, EITHER EXPRESSED OR IMPLIED, WITH RESPECT TO THIS MODEL  |
*|OR ITS FITNESS FOR A PARTICULAR PURPOSE IS CLAIMED BY TEXAS INSTRUMENTS |
*|OR THE AUTHOR.  THE MODEL IS LICENSED SOLELY ON AN "AS IS" BASIS.  THE  |
*|ENTIRE RISK AS TO ITS QUALITY AND PERFORMANCE IS WITH THE CUSTOMER.     |
* ------------------------------------------------------------------------
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TL082_0     1 2 3 4 5
*
C1   11 12 3.498E-12
C2    6  7 15.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 4.715E6 -5E6 5E6 5E6 -5E6
GA    6  0 11 12 282.8E-6
GCM   0  6 10 99 8.942E-9
ISS   3 10 DC 195.0E-6
HLIM 90  0 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100.0E3
RD1   4 11 3.536E3
RD2   4 12 3.536E3
RO1   8  5 150
RO2   7 99 150
RP    3  4 2.143E3
RSS  10 99 1.026E6
VB    9  0 DC 0
VC    3 53 DC 2.200
VE   54  4 DC 2.200
VLIM  7  8 DC 0
VLP  91  0 DC 25
VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=15.00E-12 BETA=270.1E-6 VTO=-1)
.ENDS


* MPY634_BEHAVIORAL
*****************************************************************************
* (C) COPYRIGHT 2011 TEXAS INSTRUMENTS INCORPORATED. ALL RIGHTS RESERVED.
*****************************************************************************
** THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.
** TI AND ITS LICENSORS AND SUPPLIERS MAKE NO WARRANTIES, EITHER EXPRESSED
** OR IMPLIED, WITH RESPECT TO THIS MODEL, INCLUDING THE WARRANTIES OF
** MERCHANTABILITY OR FITNESS FOR A PARTICULAR PURPOSE.  THE MODEL IS
** PROVIDED SOLELY ON AN "AS IS" BASIS.  THE ENTIRE RISK AS TO ITS QUALITY
** AND PERFORMANCE IS WITH THE CUSTOMER.
*****************************************************************************
*
* THIS MODEL IS SUBJECT TO CHANGE WITHOUT NOTICE. TEXAS INSTRUMENTS
* INCORPORATED IS NOT RESPONSIBLE FOR UPDATING THIS MODEL.
*
*****************************************************************************
*
** RELEASED BY: ANALOG ELAB DESIGN CENTER, TEXAS INSTRUMENTS INC.
* PART: MPY634
* DATE: 31JUL2011
* MODEL TYPE: BEHAVIORAL
* SIMULATOR: TINA
* SIMULATOR VERSION: 9.1.30.94 SF -TI
* EVM ORDER NUMBER: N/A
* EVM USERS GUIDE: N/A
* DATASHEET: SBFS017A � DECEMBER 1995 � REVISED DECEMBER 2004
*
* MODEL VERSION: 1.0
*
*****************************************************************************
*
* UPDATES:
*
* VERSION 1.0
*
*****************************************************************************
* THE CIRCUIT BELOW MODELS THE BEHAVIOR OF THE MPY634 FOUR QUADRANT
* MULTIPLIER BY IMPLEMENTING THE FOLLOWING TRANSFER FUNCTION:
*
*            [(X1 - X2)*(Y1 - Y2)             ]
* VOUT = A * [-------------------  - (Z1 - Z2)]
*            [         SF                     ]
*
* THE SUPPLY PINS +VS & -VS ONLY ARE USED TO CLAMP THE OUTPUT VOLTAGE TO {-VS,+VS}
* THE SCALE FACTOR OR SF HAS TO BE PROVIDED AS A DC VOLTAGE TO THE MODEL
* THE VOLTAGE AT THE SF PIN CAN IS CLAMPED INTERNALLY TO {3,10} AND MAPPED TO {0.1,10}
* THE MODEL WAS CREATED ASSUMING A SUPPLY VOLTAGE OF +/- 15 V

.SUBCKT MPY634_BEHAVIORAL_0  X1 X2 SF Y1 Y2 +VS OUT Z1 Z2 -VS

ECS3        2 0 VALUE = {LIMIT(V(SF,0),3,10)}
ECS1        3 0 VALUE = {((V(4,0)*V(5,0))/V(VF1,0)-V(6,0))*17783}
ECS4        OUT 0 VALUE = {LIMIT(V(3,0),V(-VS,0),V(+VS,0))}
ECS2        VF1 0 VALUE = {V(2,0)*9.9/7-29/7}
EZ          6 0 Z1 Z2  1
EY          5 0 Y1 Y2  1
EX          4 0 X1 X2  1

.ENDS MPY634_BEHAVIORAL_0


.END
